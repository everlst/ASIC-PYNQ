module fc_top_ip (
  input  wire        clk_i,
  input  wire        rst_n_i,
  input  wire        start_i,
  output reg         done_o,

  // === �ⲿ����RAM�ӿڣ��ӿ��Ƶ�Ԫ�ṩ�� ===
  output wire [1:0]  in_addr_o,
  input  wire [1023:0] in_data_i,

  // === ԭ��������� ===
  output wire [7:0]  final_out_wdata,
  output wire [7:0]  fc_out,
  output wire        fc_out_en,

  // === �����м���� ===
  output wire [7:0]  fc1_out_data,
  output wire        fc1_out_valid,
  output wire [7:0]  fc2_out_data,
  output wire        fc2_out_valid,
  output wire [7:0]  fc3_out_data,
  output wire        fc3_out_valid
);
  // === ԭ���źţ������� ===
  wire [   1:0] in_addr;
  wire [   9:0] w_addr;
  wire [   6:0] b_addr;

  wire [1023:0] in_data;  // t4
  wire [1023:0] w_data;  // t4
  wire [   7:0] b_data;  // t4

  wire [1023:0] mul_a;   // fc_1 �ĳ�������
  wire [1023:0] mul_b;
  wire [2047:0] mul_p;   // fc_1 �ĳ˷������2048λ��

  wire          out_wren;
  wire [  7:0] out_wdata;
  wire [   6:0] out_waddr;

  // === round_cnt ���� ===
  reg  [   7:0] round_cnt;
  always @(posedge clk_i or negedge rst_n_i) begin
    if (!rst_n_i) round_cnt <= 0;
    else if (done_o) begin
      if (round_cnt <= 8'd41) begin
        round_cnt <= round_cnt + 1'b1;
      end
    end
  end
  localparam INPUT_BLOCK_SIZE = 4;


  // start �������ݣ�����������
  wire start;
  assign start = start_i; // �ö��� start_i ���� FSM

  // ---------- RAM IP (����/Ȩ��/ƫ��) ----------

  weight_ram_rd3 u_weight_ram (
    .clka (clk_i),
    .addra(w_addr),
    .douta(w_data)
  );
  bias_ram_rd3 u_bias_ram (
    .clka (clk_i),
    .addra(b_addr),
    .douta(b_data)
  );
  // �����ⲿ���Ƶ�Ԫ����������
  assign in_data = in_data_i;
  assign in_addr_o = in_addr;
  // === ��һ�� FC (���ֽӿ�) ===
  wire done_o_1;
  fc_1 u_fc_1 (
    .clk_i  (clk_i),
    .rst_n_i(rst_n_i),
    .start_i(start),
    .done_o (done_o_1),

    .input_data_addr_o(in_addr),
    .input_data_i     (in_data),

    .weight_addr_o(w_addr),
    .weight_i     (w_data),

    .bias_addr_o(b_addr),
    .bias_i     (b_data),

    .mul_data1_o (mul_a),
    .mul_data2_o (mul_b),
    .mul_result_i(mul_p),

    .fc_output_wren_o(out_wren),
    .fc_output_data_o(out_wdata),
    .fc_output_addr_o(out_waddr)
  );

  // === ��һ�����д�� output_mem�����֣� ===
  reg [7:0] output_mem[0:127];
  always @(posedge clk_i) if (out_wren) output_mem[out_waddr] <= out_wdata[7:0];

  // === �ڶ����źţ������� ===
  wire          done_o_2;
  wire [   4:0] w_addr_2;
  wire [   4:0] b_addr_2;

  wire [1023:0] in_data_2;  // ��� output_mem -> vector
  wire [1023:0] w_data_2;
  wire [   7:0] b_data_2;

  wire [1023:0] mul_a_2;
  wire [1023:0] mul_b_2;
  wire [2047:0] mul_p_2;

  wire          out_wren_2;
  wire [  7:0] out_wdata_2;
  wire [   4:0] out_waddr_2;

  genvar j;
  generate
    for (j = 0; j < 128; j = j + 1) begin : INPUT_TO_VECTOR
      // ���ֽ�չ����ע�� index ˳����ԭʼ����һ��
      assign in_data_2[1023-8*j:1016-8*j] = output_mem[j];
    end
  endgenerate

  weight_ram_fc2 u_weight_ram_fc2 (
    .clka (clk_i),
    .addra(w_addr_2),
    .douta(w_data_2)
  );
  bias_ram_fc2 u_bias_ram_fc2 (
    .clka (clk_i),
    .addra(b_addr_2),
    .douta(b_data_2)
  );

  fc_2 u_fc_2 (
    .clk_i           (clk_i),
    .rst_n_i         (rst_n_i),
    .start_i         (done_o_1),
    .done_o          (done_o_2),
    .input_data_i    (in_data_2),
    .weight_addr_o   (w_addr_2),
    .weight_i        (w_data_2),
    .bias_addr_o     (b_addr_2),
    .bias_i          (b_data_2),
    .mul_data1_o     (mul_a_2),
    .mul_data2_o     (mul_b_2),
    .mul_result_i    (mul_p_2),
    .fc_output_wren_o(out_wren_2),
    .fc_output_data_o(out_wdata_2),
    .fc_output_addr_o(out_waddr_2)
  );

  reg [7:0] output_mem_2[0:31];
  always @(posedge clk_i) if (out_wren_2) output_mem_2[out_waddr_2] <= out_wdata_2[7:0];

  // === �������źţ������� ===
  wire          done_o_3;
  wire          w_addr_3;
  wire          b_addr_3;

  wire [ 255:0] in_data_3;
  wire [ 255:0] w_data_3;
  wire [   7:0] b_data_3;

  wire [ 255:0] mul_a_3;
  wire [ 255:0] mul_b_3;
  wire [511:0]  mul_p_3;  // ԭ��Ϊ 512 λ�����ﱣ��ԭʼλ��

  wire          out_wren_3;
  wire [  7:0] out_wdata_3;
  wire          out_waddr_3;

  generate
    for (j = 0; j < 32; j = j + 1) begin : INPUT_TO_VECTOR2
      assign in_data_3[255-8*j:248-8*j] = output_mem_2[j];
    end
  endgenerate

  weight_ram_fc3 u_weight_ram_fc3 (
    .clka (clk_i),
    .addra(w_addr_3),
    .douta(w_data_3)
  );
  bias_weight_fc3 u_bias_ram_fc3 (
    .clka (clk_i),
    .addra(b_addr_3),
    .douta(b_data_3)
  );

  fc_3 u_fc_3 (
    .clk_i           (clk_i),
    .rst_n_i         (rst_n_i),
    .start_i         (done_o_2),
    .done_o          (done_o_3),
    .input_data_i    (in_data_3),
    .weight_addr_o   (w_addr_3),
    .weight_i        (w_data_3),
    .bias_addr_o     (b_addr_3),
    .bias_i          (b_data_3),
    .mul_data1_o     (mul_a_3),
    .mul_data2_o     (mul_b_3),
    .mul_result_i    (mul_p_3),
    .fc_output_wren_o(out_wren_3),
    .fc_output_data_o(out_wdata_3),
    .fc_output_addr_o(out_waddr_3)
  );

  // �����������
  assign fc1_out_data  = out_wdata[7:0];
  assign fc1_out_valid = out_wren;
  assign fc2_out_data  = out_wdata_2[7:0];
  assign fc2_out_valid = out_wren_2;
  assign fc3_out_data  = out_wdata_3[7:0];
  assign fc3_out_valid = out_wren_3;

  assign final_out_wdata = out_wdata_3;
  assign fc_out_en = out_wren_3;
  assign fc_out    = out_wdata_3;
  always @(posedge clk_i or negedge rst_n_i) begin
    if (!rst_n_i) done_o <= 0;
    else  begin
      done_o     = done_o_3;
    end
  end

  // ===================================================
  // ========== ����˷��� + FSM �����߼� ================
  // ===================================================
  // ����ʹ��һ�� NUM_MULTIPLIERS = 128 �� multiplier_array ��Ϊ����˷���
  // mul_a_shared/mul_b_shared ���Ϊ 1024 (��ԭ 128 ������������һ��)
  // mul_p_shared ���Ϊ 2048 (��ԭ 128 �����������һ��)
  // fc_1 / fc_2 �ڴ� 2048 λ��� -> ֱ��ʹ�� mul_p_shared
  // fc_3 �ڴ���С�Ľ�� (512 λ) -> ʹ�� mul_p_shared[511:0] ��Ϊ������

  // FSM ״̬����
  localparam S_IDLE = 2'd0,
             S_FC1  = 2'd1,
             S_FC2  = 2'd2,
             S_FC3  = 2'd3;

  reg [1:0] fc_state, fc_state_next;

  // ״̬�Ĵ�
  always @(posedge clk_i or negedge rst_n_i) begin
    if (!rst_n_i) fc_state <= S_IDLE;
    else fc_state <= fc_state_next;
  end

  // ��һ״̬����߼�������ʹ�ø��� done �źţ�
  always @(*) begin
    fc_state_next = fc_state;
    case (fc_state)
      S_IDLE: begin
        if (start) fc_state_next = S_FC1;
        else fc_state_next = S_IDLE;
      end
      S_FC1: begin
        if (done_o_1) fc_state_next = S_FC2;
        else fc_state_next = S_FC1;
      end
      S_FC2: begin
        if (done_o_2) fc_state_next = S_FC3;
        else fc_state_next = S_FC2;
      end
      S_FC3: begin
        if (done_o_3) fc_state_next = S_IDLE;
        else fc_state_next = S_FC3;
      end
      default: fc_state_next = S_IDLE;
    endcase
  end

  // ����˷��������루1024 λ each��
  reg  [1023:0] mul_a_shared;
  reg  [1023:0] mul_b_shared;
  wire [2047:0] mul_p_shared;

  // ���ݵ�ǰ״̬�Ѷ�Ӧ��� mul_a_x/mul_b_x ���빲��˷���
  // �Խ�խ�ĵ���������������չ�� 1024 λ
  always @(*) begin
    case (fc_state)
      S_FC1: begin
        mul_a_shared = mul_a;     // fc_1 ԭʼ 1024 λ����
        mul_b_shared = mul_b;
      end
      S_FC2: begin
        mul_a_shared = mul_a_2;   // fc_2 ԭʼ 1024 λ����
        mul_b_shared = mul_b_2;
      end
      S_FC3: begin
        // fc_3 ֻ�� 256 λ���� (mul_a_3 / mul_b_3)
        // ����λ�ŵ� shared �ĵ� 256 λ�� ��λ�� 0
        mul_a_shared = {768'd0, mul_a_3};
        mul_b_shared = {768'd0, mul_b_3};
      end
      default: begin
        mul_a_shared = 1024'd0;
        mul_b_shared = 1024'd0;
      end
    endcase
  end

  // ����˷���ʵ������һ����
  multiplier_array #(
    .NUM_MULTIPLIERS(128)
  ) u_mult_array_shared (
    .clk_i(clk_i),
    .mul_a(mul_a_shared),
    .mul_b(mul_b_shared),
    .mul_p(mul_p_shared)
  );

  // ������˷�������ַ��ظ���� mul_result �ӿ�
  // fc_1 �� fc_2 ��Ҫ������ 2048 λ���
  // fc_3 ������С�Ľ����ȡ��λ���֣�512 λ��
  // ע�⣺ԭ�� fc_3 mul_p_3 ���д�� [512:0] (513 bits)��Ϊ�˼������������Ϊ 513 λ����λ��
  // ���ԭʼ fc_3 ��ʹ�� 512 λ������Ӧ������ģ��
  assign mul_p  = mul_p_shared;              // 2048 λ -> fc_1
  assign mul_p_2 = mul_p_shared;             // 2048 λ -> fc_2
  
  // �ѵ� 512 λ�� fc_3��ԭ�ȶ��� mul_p_3 �� [512:0]��
  // ������ fc_3 ʵ�ʽ��� 512 λ����������������Ϊ [511:0]
  assign mul_p_3 =  mul_p_shared[511:0]; // ��λ padding 0 -> �ܿ�� 513 λ

  // ===================================================
  // End of shared multiplier + FSM
  // ===================================================

endmodule

